module 32bit_MUL();
endmodule
