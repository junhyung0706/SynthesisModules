module 1bit_HA();
endmodule
