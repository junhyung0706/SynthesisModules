module Top();
endmodule
