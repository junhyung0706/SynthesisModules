module 1bit_FA();
endmodule
