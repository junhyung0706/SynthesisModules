module 32bit_RCA();
endmodule
