module 32bit_MUL(
input [31:0] A,
input [7:0] B,
output [39:0] Y
);

wire [15:0] w1,w2,w3;

//              a&b,       Sin, Cin, Sout, Cout
1bit_FA FA0_0(A[0] & B[0], 1'b0, 1'b0, Y[0], w1[1]); //A[0]*B[0]을 수행하는 FA
1bit_FA FA0_1(A[0] & B[1], 1'b0, 1'b0, w1[2], w1[3]); //A[0]*B[1]을 수행하는 FA
1bit_FA FA0_2(A[0] & B[2], 1'b0, 1'b0, w1[4], w1[5]);
1bit_FA FA0_3(A[0] & B[3], 1'b0, 1'b0, w1[6], w1[7]);
1bit_FA FA0_4(A[0] & B[4], 1'b0, 1'b0, w1[8], w1[9]);
1bit_FA FA0_5(A[0] & B[5], 1'b0, 1'b0, w1[10], w1[11]);
1bit_FA FA0_6(A[0] & B[6], 1'b0, 1'b0, w1[12], w1[13]);
1bit_FA FA0_7(A[0] & B[7], 1'b0, 1'b0, w1[14], w1[15]);

1bit_FA FA1_0(A[1]& B[0], w1[2], w1[1], Y[1], w2[1]);
1bit_FA FA1_1(A[1]& B[1], w1[4], w1[3], w2[2], w2[3]);
1bit_FA FA1_2(A[1]& B[2], w1[6], w1[5], w2[4], w2[5]);
1bit_FA FA1_3(A[1]& B[3], w1[8] ,w1[7], w2[6], w2[7]);
1bit_FA FA1_4(A[1]& B[4], w1[10], w1[9], w2[8], w2[9]);
1bit_FA FA1_5(A[1]& B[5], w1[12], w1[11], w2[10], w2[11]);
1bit_FA FA1_6(A[1]& B[6], w1[14], w1[13], w2[12], w2[13]);
1bit_FA FA1_7(A[1]& B[7], 1'b0, w1[14], w2[14], w2[15]);

1bit_FA FA2_0(A[2]& B[0], w2[2], w2[1], Y[2], w3[1]);
1bit_FA FA2_1(A[2]& B[1], w2[4], w2[3], w3[2], w3[3]);
1bit_FA FA2_2(A[2]& B[2], w2[6], w2[5], w3[4], w3[5]);
1bit_FA FA2_3(A[2]& B[3], w2[8], w2[7], w3[6], w3[7]);
1bit_FA FA2_4(A[2]& B[4], w2[10], w2[9], w3[8], w3[9]);
1bit_FA FA2_5(A[2]& B[5], w2[12], w2[11], w3[10], w3[11]);
1bit_FA FA2_6(A[2]& B[6], w2[14], w2[13], w3[12], w3[13]);
1bit_FA FA2_7(A[2]& B[7], 1'b0, w2[14], w3[14], w3[15]);




endmodule