module 32bit_CSA();
endmodule
