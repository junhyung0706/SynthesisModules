module bit32_MUL(
input [31:0] A,
input [7:0] B,
output [39:0] Y
);

wire [14:0] w1,w2,w3,w4,w5,w6,w7,w8,w9,w10;
wire [14:0] w11,w12,w13,w14,w15,w16,w17,w18,w19,w20;
wire [14:0] w21,w22,w23,w24,w25,w26,w27,w28,w29,w30,w31,w32;
wire [7:0] LastCarry;

//              a&b,       Sin, Cin, Sout, Cout
bit1_FA FA0_0(A[0] & B[0], 1'b0, 1'b0, Y[0], w1[0]); //A[0]*B[0]을 수행하는 FA
bit1_FA FA0_1(A[0] & B[1], 1'b0, 1'b0, w1[1], w1[2]); //A[0]*B[1]을 수행하는 FA
bit1_FA FA0_2(A[0] & B[2], 1'b0, 1'b0, w1[3], w1[4]);
bit1_FA FA0_3(A[0] & B[3], 1'b0, 1'b0, w1[5], w1[6]);
bit1_FA FA0_4(A[0] & B[4], 1'b0, 1'b0, w1[7], w1[8]);
bit1_FA FA0_5(A[0] & B[5], 1'b0, 1'b0, w1[9], w1[10]);
bit1_FA FA0_6(A[0] & B[6], 1'b0, 1'b0, w1[11], w1[12]);
bit1_FA FA0_7(A[0] & B[7], 1'b0, 1'b0, w1[13], w1[14]);

bit1_FA FA1_0(A[1]& B[0], w1[1], w1[0], Y[1], w2[0]);
bit1_FA FA1_1(A[1]& B[1], w1[3], w1[2], w2[1], w2[2]);
bit1_FA FA1_2(A[1]& B[2], w1[5], w1[4], w2[3], w2[4]);
bit1_FA FA1_3(A[1]& B[3], w1[7] ,w1[6], w2[5], w2[6]);
bit1_FA FA1_4(A[1]& B[4], w1[9], w1[8], w2[7], w2[8]);
bit1_FA FA1_5(A[1]& B[5], w1[11], w1[10], w2[9], w2[10]);
bit1_FA FA1_6(A[1]& B[6], w1[13], w1[12], w2[11], w2[12]);
bit1_FA FA1_7(A[1]& B[7], 1'b0, w1[14], w2[13], w2[14]);

bit1_FA FA2_0(A[2]& B[0], w2[1], w2[0], Y[2], w3[0]);
bit1_FA FA2_1(A[2]& B[1], w2[3], w2[2], w3[1], w3[2]);
bit1_FA FA2_2(A[2]& B[2], w2[5], w2[4], w3[3], w3[4]);
bit1_FA FA2_3(A[2]& B[3], w2[7], w2[6], w3[5], w3[6]);
bit1_FA FA2_4(A[2]& B[4], w2[9], w2[8], w3[7], w3[8]);
bit1_FA FA2_5(A[2]& B[5], w2[11], w2[10], w3[9], w3[10]);
bit1_FA FA2_6(A[2]& B[6], w2[13], w2[12], w3[11], w3[12]);
bit1_FA FA2_7(A[2]& B[7], 1'b0, w2[14], w3[13], w3[14]);

bit1_FA FA3_0(A[3]& B[0], w3[1], w3[0], Y[3], w4[0]);
bit1_FA FA3_1(A[3]& B[1], w3[3], w3[2], w4[1], w4[2]);
bit1_FA FA3_2(A[3]& B[2], w3[5], w3[4], w4[3], w4[4]);
bit1_FA FA3_3(A[3]& B[3], w3[7], w3[6], w4[5], w4[6]);
bit1_FA FA3_4(A[3]& B[4], w3[9], w3[8], w4[7], w4[8]);
bit1_FA FA3_5(A[3]& B[5], w3[11], w3[10], w4[9], w4[10]);
bit1_FA FA3_6(A[3]& B[6], w3[13], w3[12], w4[11], w4[12]);
bit1_FA FA3_7(A[3]& B[7], 1'b0, w3[14], w4[13], w4[14]);

bit1_FA FA4_0(A[4]& B[0], w4[1], w4[0], Y[4], w5[0]);
bit1_FA FA4_1(A[4]& B[1], w4[3], w4[2], w5[1], w5[2]);
bit1_FA FA4_2(A[4]& B[2], w4[5], w4[4], w5[3], w5[4]);
bit1_FA FA4_3(A[4]& B[3], w4[7], w4[6], w5[5], w5[6]);
bit1_FA FA4_4(A[4]& B[4], w4[9], w4[8], w5[7], w5[8]);
bit1_FA FA4_5(A[4]& B[5], w4[11], w4[10], w5[9], w5[10]);
bit1_FA FA4_6(A[4]& B[6], w4[13], w4[12], w5[11], w5[12]);
bit1_FA FA4_7(A[4]& B[7], 1'b0, w4[14], w5[13], w5[14]);

bit1_FA FA5_0(A[5]& B[0], w5[1], w5[0], Y[5], w6[0]);
bit1_FA FA5_1(A[5]& B[1], w5[3], w5[2], w6[1], w6[2]);
bit1_FA FA5_2(A[5]& B[2], w5[5], w5[4], w6[3], w6[4]);
bit1_FA FA5_3(A[5]& B[3], w5[7], w5[6], w6[5], w6[6]);
bit1_FA FA5_4(A[5]& B[4], w5[9], w5[8], w6[7], w6[8]);
bit1_FA FA5_5(A[5]& B[5], w5[11], w5[10], w6[9], w6[10]);
bit1_FA FA5_6(A[5]& B[6], w5[13], w5[12], w6[11], w6[12]);
bit1_FA FA5_7(A[5]& B[7], 1'b0, w5[14], w6[13], w6[14]);

bit1_FA FA6_0(A[6]& B[0], w6[1], w6[0], Y[6], w7[0]);
bit1_FA FA6_1(A[6]& B[1], w6[3], w6[2], w7[1], w7[2]);
bit1_FA FA6_2(A[6]& B[2], w6[5], w6[4], w7[3], w7[4]);
bit1_FA FA6_3(A[6]& B[3], w6[7], w6[6], w7[5], w7[6]);
bit1_FA FA6_4(A[6]& B[4], w6[9], w6[8], w7[7], w7[8]);
bit1_FA FA6_5(A[6]& B[5], w6[11], w6[10], w7[9], w7[10]);
bit1_FA FA6_6(A[6]& B[6], w6[13], w6[12], w7[11], w7[12]);
bit1_FA FA6_7(A[6]& B[7], 1'b0, w6[14], w7[13], w7[14]);

bit1_FA FA7_0(A[7]& B[0], w7[1], w7[0], Y[7], w8[0]);
bit1_FA FA7_1(A[7]& B[1], w7[3], w7[2], w8[1], w8[2]);
bit1_FA FA7_2(A[7]& B[2], w7[5], w7[4], w8[3], w8[4]);
bit1_FA FA7_3(A[7]& B[3], w7[7], w7[6], w8[5], w8[6]);
bit1_FA FA7_4(A[7]& B[4], w7[9], w7[8], w8[7], w8[8]);
bit1_FA FA7_5(A[7]& B[5], w7[11], w7[10], w8[9], w8[10]);
bit1_FA FA7_6(A[7]& B[6], w7[13], w7[12], w8[11], w8[12]);
bit1_FA FA7_7(A[7]& B[7], 1'b0, w7[14], w8[13], w8[14]);

bit1_FA FA8_0(A[8]& B[0], w8[1], w8[0], Y[8], w9[0]);
bit1_FA FA8_1(A[8]& B[1], w8[3], w8[2], w9[1], w9[2]);
bit1_FA FA8_2(A[8]& B[2], w8[5], w8[4], w9[3], w9[4]);
bit1_FA FA8_3(A[8]& B[3], w8[7], w8[6], w9[5], w9[6]);
bit1_FA FA8_4(A[8]& B[4], w8[9], w8[8], w9[7], w9[8]);
bit1_FA FA8_5(A[8]& B[5], w8[11], w8[10], w9[9], w9[10]);
bit1_FA FA8_6(A[8]& B[6], w8[13], w8[12], w9[11], w9[12]);
bit1_FA FA8_7(A[8]& B[7], 1'b0, w8[14], w9[13], w9[14]);

bit1_FA FA9_0(A[9]& B[0], w9[1], w9[0], Y[9], w10[0]);
bit1_FA FA9_1(A[9]& B[1], w9[3], w9[2], w10[1], w10[2]);
bit1_FA FA9_2(A[9]& B[2], w9[5], w9[4], w10[3], w10[4]);
bit1_FA FA9_3(A[9]& B[3], w9[7], w9[6], w10[5], w10[6]);
bit1_FA FA9_4(A[9]& B[4], w9[9], w9[8], w10[7], w10[8]);
bit1_FA FA9_5(A[9]& B[5], w9[11], w9[10], w10[9], w10[10]);
bit1_FA FA9_6(A[9]& B[6], w9[13], w9[12], w10[11], w10[12]);
bit1_FA FA9_7(A[9]& B[7], 1'b0, w9[14], w10[13], w10[14]);

bit1_FA FA10_0(A[10]& B[0], w10[1], w10[0], Y[10], w11[0]);
bit1_FA FA10_1(A[10]& B[1], w10[3], w10[2], w11[1], w11[2]);
bit1_FA FA10_2(A[10]& B[2], w10[5], w10[4], w11[3], w11[4]);
bit1_FA FA10_3(A[10]& B[3], w10[7], w10[6], w11[5], w11[6]);
bit1_FA FA10_4(A[10]& B[4], w10[9], w10[8], w11[7], w11[8]);
bit1_FA FA10_5(A[10]& B[5], w10[11], w10[10], w11[9], w11[10]);
bit1_FA FA10_6(A[10]& B[6], w10[13], w10[12], w11[11], w11[12]);
bit1_FA FA10_7(A[10]& B[7], 1'b0, w10[14], w11[13], w11[14]);

bit1_FA FA11_0(A[11]& B[0], w11[1], w11[0], Y[11], w12[0]);
bit1_FA FA11_1(A[11]& B[1], w11[3], w11[2], w12[1], w12[2]);
bit1_FA FA11_2(A[11]& B[2], w11[5], w11[4], w12[3], w12[4]);
bit1_FA FA11_3(A[11]& B[3], w11[7], w11[6], w12[5], w12[6]);
bit1_FA FA11_4(A[11]& B[4], w11[9], w11[8], w12[7], w12[8]);
bit1_FA FA11_5(A[11]& B[5], w11[11], w11[10], w12[9], w12[10]);
bit1_FA FA11_6(A[11]& B[6], w11[13], w11[12], w12[11], w12[12]);
bit1_FA FA11_7(A[11]& B[7], 1'b0, w11[14], w12[13], w12[14]);

bit1_FA FA12_0(A[12]& B[0], w12[1], w12[0], Y[12], w13[0]);
bit1_FA FA12_1(A[12]& B[1], w12[3], w12[2], w13[1], w13[2]);
bit1_FA FA12_2(A[12]& B[2], w12[5], w12[4], w13[3], w13[4]);
bit1_FA FA12_3(A[12]& B[3], w12[7], w12[6], w13[5], w13[6]);
bit1_FA FA12_4(A[12]& B[4], w12[9], w12[8], w13[7], w13[8]);
bit1_FA FA12_5(A[12]& B[5], w12[11], w12[10], w13[9], w13[10]);
bit1_FA FA12_6(A[12]& B[6], w12[13], w12[12], w13[11], w13[12]);
bit1_FA FA12_7(A[12]& B[7], 1'b0, w12[14], w13[13], w13[14]);

bit1_FA FA13_0(A[13]& B[0], w13[1], w13[0], Y[13], w14[0]);
bit1_FA FA13_1(A[13]& B[1], w13[3], w13[2], w14[1], w14[2]);
bit1_FA FA13_2(A[13]& B[2], w13[5], w13[4], w14[3], w14[4]);
bit1_FA FA13_3(A[13]& B[3], w13[7], w13[6], w14[5], w14[6]);
bit1_FA FA13_4(A[13]& B[4], w13[9], w13[8], w14[7], w14[8]);
bit1_FA FA13_5(A[13]& B[5], w13[11], w13[10], w14[9], w14[10]);
bit1_FA FA13_6(A[13]& B[6], w13[13], w13[12], w14[11], w14[12]);
bit1_FA FA13_7(A[13]& B[7], 1'b0, w13[14], w14[13], w14[14]);

bit1_FA FA14_0(A[14]& B[0], w14[1], w14[0], Y[14], w15[0]);
bit1_FA FA14_1(A[14]& B[1], w14[3], w14[2], w15[1], w15[2]);
bit1_FA FA14_2(A[14]& B[2], w14[5], w14[4], w15[3], w15[4]);
bit1_FA FA14_3(A[14]& B[3], w14[7], w14[6], w15[5], w15[6]);
bit1_FA FA14_4(A[14]& B[4], w14[9], w14[8], w15[7], w15[8]);
bit1_FA FA14_5(A[14]& B[5], w14[11], w14[10], w15[9], w15[10]);
bit1_FA FA14_6(A[14]& B[6], w14[13], w14[12], w15[11], w15[12]);
bit1_FA FA14_7(A[14]& B[7], 1'b0, w14[14], w15[13], w15[14]);

bit1_FA FA15_0(A[15]& B[0], w15[1], w15[0], Y[15], w16[0]);
bit1_FA FA15_1(A[15]& B[1], w15[3], w15[2], w16[1], w16[2]);
bit1_FA FA15_2(A[15]& B[2], w15[5], w15[4], w16[3], w16[4]);
bit1_FA FA15_3(A[15]& B[3], w15[7], w15[6], w16[5], w16[6]);
bit1_FA FA15_4(A[15]& B[4], w15[9], w15[8], w16[7], w16[8]);
bit1_FA FA15_5(A[15]& B[5], w15[11], w15[10], w16[9], w16[10]);
bit1_FA FA15_6(A[15]& B[6], w15[13], w15[12], w16[11], w16[12]);
bit1_FA FA15_7(A[15]& B[7], 1'b0, w15[14], w16[13], w16[14]);

bit1_FA FA16_0(A[16]& B[0], w16[1], w16[0], Y[16], w17[0]);
bit1_FA FA16_1(A[16]& B[1], w16[3], w16[2], w17[1], w17[2]);
bit1_FA FA16_2(A[16]& B[2], w16[5], w16[4], w17[3], w17[4]);
bit1_FA FA16_3(A[16]& B[3], w16[7], w16[6], w17[5], w17[6]);
bit1_FA FA16_4(A[16]& B[4], w16[9], w16[8], w17[7], w17[8]);
bit1_FA FA16_5(A[16]& B[5], w16[11], w16[10], w17[9], w17[10]);
bit1_FA FA16_6(A[16]& B[6], w16[13], w16[12], w17[11], w17[12]);
bit1_FA FA16_7(A[16]& B[7], 1'b0, w16[14], w17[13], w17[14]);

bit1_FA FA17_0(A[17]& B[0], w17[1], w17[0], Y[17], w18[0]);
bit1_FA FA17_1(A[17]& B[1], w17[3], w17[2], w18[1], w18[2]);
bit1_FA FA17_2(A[17]& B[2], w17[5], w17[4], w18[3], w18[4]);
bit1_FA FA17_3(A[17]& B[3], w17[7], w17[6], w18[5], w18[6]);
bit1_FA FA17_4(A[17]& B[4], w17[9], w17[8], w18[7], w18[8]);
bit1_FA FA17_5(A[17]& B[5], w17[11], w17[10], w18[9], w18[10]);
bit1_FA FA17_6(A[17]& B[6], w17[13], w17[12], w18[11], w18[12]);
bit1_FA FA17_7(A[17]& B[7], 1'b0, w17[14], w18[13], w18[14]);

bit1_FA FA18_0(A[18]& B[0], w18[1], w18[0], Y[18], w19[0]);
bit1_FA FA18_1(A[18]& B[1], w18[3], w18[2], w19[1], w19[2]);
bit1_FA FA18_2(A[18]& B[2], w18[5], w18[4], w19[3], w19[4]);
bit1_FA FA18_3(A[18]& B[3], w18[7], w18[6], w19[5], w19[6]);
bit1_FA FA18_4(A[18]& B[4], w18[9], w18[8], w19[7], w19[8]);
bit1_FA FA18_5(A[18]& B[5], w18[11], w18[10], w19[9], w19[10]);
bit1_FA FA18_6(A[18]& B[6], w18[13], w18[12], w19[11], w19[12]);
bit1_FA FA18_7(A[18]& B[7], 1'b0, w18[14], w19[13], w19[14]);

bit1_FA FA19_0(A[19]& B[0], w19[1], w19[0], Y[19], w20[0]);
bit1_FA FA19_1(A[19]& B[1], w19[3], w19[2], w20[1], w20[2]);
bit1_FA FA19_2(A[19]& B[2], w19[5], w19[4], w20[3], w20[4]);
bit1_FA FA19_3(A[19]& B[3], w19[7], w19[6], w20[5], w20[6]);
bit1_FA FA19_4(A[19]& B[4], w19[9], w19[8], w20[7], w20[8]);
bit1_FA FA19_5(A[19]& B[5], w19[11], w19[10], w20[9], w20[10]);
bit1_FA FA19_6(A[19]& B[6], w19[13], w19[12], w20[11], w20[12]);
bit1_FA FA19_7(A[19]& B[7], 1'b0, w19[14], w20[13], w20[14]);

bit1_FA FA20_0(A[20]& B[0], w20[1], w20[0], Y[20], w21[0]);
bit1_FA FA20_1(A[20]& B[1], w20[3], w20[2], w21[1], w21[2]);
bit1_FA FA20_2(A[20]& B[2], w20[5], w20[4], w21[3], w21[4]);
bit1_FA FA20_3(A[20]& B[3], w20[7], w20[6], w21[5], w21[6]);
bit1_FA FA20_4(A[20]& B[4], w20[9], w20[8], w21[7], w21[8]);
bit1_FA FA20_5(A[20]& B[5], w20[11], w20[10], w21[9], w21[10]);
bit1_FA FA20_6(A[20]& B[6], w20[13], w20[12], w21[11], w21[12]);
bit1_FA FA20_7(A[20]& B[7], 1'b0, w20[14], w21[13], w21[14]);

bit1_FA FA21_0(A[21]& B[0], w21[1], w21[0], Y[21], w22[0]);
bit1_FA FA21_1(A[21]& B[1], w21[3], w21[2], w22[1], w22[2]);
bit1_FA FA21_2(A[21]& B[2], w21[5], w21[4], w22[3], w22[4]);
bit1_FA FA21_3(A[21]& B[3], w21[7], w21[6], w22[5], w22[6]);
bit1_FA FA21_4(A[21]& B[4], w21[9], w21[8], w22[7], w22[8]);
bit1_FA FA21_5(A[21]& B[5], w21[11], w21[10], w22[9], w22[10]);
bit1_FA FA21_6(A[21]& B[6], w21[13], w21[12], w22[11], w22[12]);
bit1_FA FA21_7(A[21]& B[7], 1'b0, w21[14], w22[13], w22[14]);

bit1_FA FA22_0(A[22]& B[0], w22[1], w22[0], Y[22], w23[0]);
bit1_FA FA22_1(A[22]& B[1], w22[3], w22[2], w23[1], w23[2]);
bit1_FA FA22_2(A[22]& B[2], w22[5], w22[4], w23[3], w23[4]);
bit1_FA FA22_3(A[22]& B[3], w22[7], w22[6], w23[5], w23[6]);
bit1_FA FA22_4(A[22]& B[4], w22[9], w22[8], w23[7], w23[8]);
bit1_FA FA22_5(A[22]& B[5], w22[11], w22[10], w23[9], w23[10]);
bit1_FA FA22_6(A[22]& B[6], w22[13], w22[12], w23[11], w23[12]);
bit1_FA FA22_7(A[22]& B[7], 1'b0, w22[14], w23[13], w23[14]);

bit1_FA FA23_0(A[23]& B[0], w23[1], w23[0], Y[23], w24[0]);
bit1_FA FA23_1(A[23]& B[1], w23[3], w23[2], w24[1], w24[2]);
bit1_FA FA23_2(A[23]& B[2], w23[5], w23[4], w24[3], w24[4]);
bit1_FA FA23_3(A[23]& B[3], w23[7], w23[6], w24[5], w24[6]);
bit1_FA FA23_4(A[23]& B[4], w23[9], w23[8], w24[7], w24[8]);
bit1_FA FA23_5(A[23]& B[5], w23[11], w23[10], w24[9], w24[10]);
bit1_FA FA23_6(A[23]& B[6], w23[13], w23[12], w24[11], w24[12]);
bit1_FA FA23_7(A[23]& B[7], 1'b0, w23[14], w24[13], w24[14]);

bit1_FA FA24_0(A[24]& B[0], w24[1], w24[0], Y[24], w25[0]);
bit1_FA FA24_1(A[24]& B[1], w24[3], w24[2], w25[1], w25[2]);
bit1_FA FA24_2(A[24]& B[2], w24[5], w24[4], w25[3], w25[4]);
bit1_FA FA24_3(A[24]& B[3], w24[7], w24[6], w25[5], w25[6]);
bit1_FA FA24_4(A[24]& B[4], w24[9], w24[8], w25[7], w25[8]);
bit1_FA FA24_5(A[24]& B[5], w24[11], w24[10], w25[9], w25[10]);
bit1_FA FA24_6(A[24]& B[6], w24[13], w24[12], w25[11], w25[12]);
bit1_FA FA24_7(A[24]& B[7], 1'b0, w24[14], w25[13], w25[14]);

bit1_FA FA25_0(A[25]& B[0], w25[1], w25[0], Y[25], w26[0]);
bit1_FA FA25_1(A[25]& B[1], w25[3], w25[2], w26[1], w26[2]);
bit1_FA FA25_2(A[25]& B[2], w25[5], w25[4], w26[3], w26[4]);
bit1_FA FA25_3(A[25]& B[3], w25[7], w25[6], w26[5], w26[6]);
bit1_FA FA25_4(A[25]& B[4], w25[9], w25[8], w26[7], w26[8]);
bit1_FA FA25_5(A[25]& B[5], w25[11], w25[10], w26[9], w26[10]);
bit1_FA FA25_6(A[25]& B[6], w25[13], w25[12], w26[11], w26[12]);
bit1_FA FA25_7(A[25]& B[7], 1'b0, w25[14], w26[13], w26[14]);

bit1_FA FA26_0(A[26]& B[0], w26[1], w26[0], Y[26], w27[0]);
bit1_FA FA26_1(A[26]& B[1], w26[3], w26[2], w27[1], w27[2]);
bit1_FA FA26_2(A[26]& B[2], w26[5], w26[4], w27[3], w27[4]);
bit1_FA FA26_3(A[26]& B[3], w26[7], w26[6], w27[5], w27[6]);
bit1_FA FA26_4(A[26]& B[4], w26[9], w26[8], w27[7], w27[8]);
bit1_FA FA26_5(A[26]& B[5], w26[11], w26[10], w27[9], w27[10]);
bit1_FA FA26_6(A[26]& B[6], w26[13], w26[12], w27[11], w27[12]);
bit1_FA FA26_7(A[26]& B[7], 1'b0, w26[14], w27[13], w27[14]);

bit1_FA FA27_0(A[27]& B[0], w27[1], w27[0], Y[27], w28[0]);
bit1_FA FA27_1(A[27]& B[1], w27[3], w27[2], w28[1], w28[2]);
bit1_FA FA27_2(A[27]& B[2], w27[5], w27[4], w28[3], w28[4]);
bit1_FA FA27_3(A[27]& B[3], w27[7], w27[6], w28[5], w28[6]);
bit1_FA FA27_4(A[27]& B[4], w27[9], w27[8], w28[7], w28[8]);
bit1_FA FA27_5(A[27]& B[5], w27[11], w27[10], w28[9], w28[10]);
bit1_FA FA27_6(A[27]& B[6], w27[13], w27[12], w28[11], w28[12]);
bit1_FA FA27_7(A[27]& B[7], 1'b0, w27[14], w28[13], w28[14]);

bit1_FA FA28_0(A[28]& B[0], w28[1], w28[0], Y[28], w29[0]);
bit1_FA FA28_1(A[28]& B[1], w28[3], w28[2], w29[1], w29[2]);
bit1_FA FA28_2(A[28]& B[2], w28[5], w28[4], w29[3], w29[4]);
bit1_FA FA28_3(A[28]& B[3], w28[7], w28[6], w29[5], w29[6]);
bit1_FA FA28_4(A[28]& B[4], w28[9], w28[8], w29[7], w29[8]);
bit1_FA FA28_5(A[28]& B[5], w28[11], w28[10], w29[9], w29[10]);
bit1_FA FA28_6(A[28]& B[6], w28[13], w28[12], w29[11], w29[12]);
bit1_FA FA28_7(A[28]& B[7], 1'b0, w28[14], w29[13], w29[14]);

bit1_FA FA29_0(A[29]& B[0], w29[1], w29[0], Y[29], w30[0]);
bit1_FA FA29_1(A[29]& B[1], w29[3], w29[2], w30[1], w30[2]);
bit1_FA FA29_2(A[29]& B[2], w29[5], w29[4], w30[3], w30[4]);
bit1_FA FA29_3(A[29]& B[3], w29[7], w29[6], w30[5], w30[6]);
bit1_FA FA29_4(A[29]& B[4], w29[9], w29[8], w30[7], w30[8]);
bit1_FA FA29_5(A[29]& B[5], w29[11], w29[10], w30[9], w30[10]);
bit1_FA FA29_6(A[29]& B[6], w29[13], w29[12], w30[11], w30[12]);
bit1_FA FA29_7(A[29]& B[7], 1'b0, w29[14], w30[13], w30[14]);

bit1_FA FA30_0(A[30]& B[0], w30[1], w30[0], Y[30], w31[0]);
bit1_FA FA30_1(A[30]& B[1], w30[3], w30[2], w31[1], w31[2]);
bit1_FA FA30_2(A[30]& B[2], w30[5], w30[4], w31[3], w31[4]);
bit1_FA FA30_3(A[30]& B[3], w30[7], w30[6], w31[5], w31[6]);
bit1_FA FA30_4(A[30]& B[4], w30[9], w30[8], w31[7], w31[8]);
bit1_FA FA30_5(A[30]& B[5], w30[11], w30[10], w31[9], w31[10]);
bit1_FA FA30_6(A[30]& B[6], w30[13], w30[12], w31[11], w31[12]);
bit1_FA FA30_7(A[30]& B[7], 1'b0, w30[14], w31[13], w31[14]);

bit1_FA FA31_0(A[31]& B[0], w31[1], w31[0], Y[31], w32[0]);
bit1_FA FA31_1(A[31]& B[1], w31[3], w31[2], w32[1], w32[2]);
bit1_FA FA31_2(A[31]& B[2], w31[5], w31[4], w32[3], w32[4]);
bit1_FA FA31_3(A[31]& B[3], w31[7], w31[6], w32[5], w32[6]);
bit1_FA FA31_4(A[31]& B[4], w31[9], w31[8], w32[7], w32[8]);
bit1_FA FA31_5(A[31]& B[5], w31[11], w31[10], w32[9], w32[10]);
bit1_FA FA31_6(A[31]& B[6], w31[13], w31[12], w32[11], w32[12]);
bit1_FA FA31_7(A[31]& B[7], 1'b0, w31[14], w32[13], w32[14]);

//마지막 줄의 모듈들
bit1_FA FA0(w32[1], w32[0], 1'b0, Y[32], LastCarry[0]);
bit1_FA FA1(w32[3], w32[2], LastCarry[0], Y[33], LastCarry[1]);
bit1_FA FA2(w32[5], w32[4], LastCarry[1], Y[34], LastCarry[2]);
bit1_FA FA3(w32[7], w32[6], LastCarry[2], Y[35], LastCarry[3]);
bit1_FA FA4(w32[9], w32[8], LastCarry[3], Y[36], LastCarry[4]);
bit1_FA FA5(w32[11], w32[10], LastCarry[4], Y[37], LastCarry[5]);
bit1_FA FA6(w32[13], w32[12], LastCarry[5], Y[38], LastCarry[6]);
bit1_FA FA7(1'b0, w32[14], LastCarry[6], Y[39], LastCarry[7]);

endmodule
