module 4bit_RCA();
endmodule
