module 32bit_MUL(
    input [31:0] A,
    input [7:0] B,
    output [39:0] Y
);


endmodule
